(*blackbox*)
module v2f_rolling_accumulate(
	input signed [31:0] A, // Accumulate
	output [31:0] Y); //Sum of data
endmodule